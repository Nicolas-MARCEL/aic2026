magic
tech sky130A
timestamp 1768757060
<< locali >>
rect -48 -200 48 76
rect 533 -200 629 3
rect -48 -296 629 -200
rect 299 -300 400 -296
<< metal1 >>
rect -92 -64 668 2064
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xo0<1>
timestamp 1740610800
transform 1 0 0 0 1 400
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xo1<0>
timestamp 1740610800
transform 1 0 0 0 1 1200
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xo1<1>
timestamp 1740610800
transform 1 0 0 0 1 1600
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xo1
timestamp 1740610800
transform 1 0 0 0 1 800
box -92 -64 668 464
<< properties >>
string FIXED_BBOX 0 0 576 2000
<< end >>
